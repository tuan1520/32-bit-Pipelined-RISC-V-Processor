module bin2bcd(
  input  logic [31:0] i_bin,
  output logic [31:0] o_bcd
);
  assign o_bcd = i_bin; // placeholder
endmodule
